module Forwarding(p0, p1, forwardP0, forwardP1);

endmodule
